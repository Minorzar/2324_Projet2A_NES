-- interrupt_and_reset_control.vhd
--
-- This VHDL module implements "Interrupt and Reset Control Logic".
--
-- Description:
--	

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity interrupt_and_reset_control is
	Port (
		i_placeholder				: in std_logic;						-- Input signal
		o_placeholder				: in std_logic;						-- Output signal
	);
end interrupt_and_reset_control;

architecture Behavioral of interrupt_and_reset_control is
	signal placeholder			: std_logic;
begin

end Behavioral;

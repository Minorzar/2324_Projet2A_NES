library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; 


entity ALU is 

end ALU; 


architecture ALU_rtf of ALU is
begin

end ALU_rft; 
-- decode_rom.vhd
-- placeholder.vhd
--
-- This VHDL module implements "Placeholder".
--
-- Description:
--	

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity placeholder is
	Port (
		i_placeholder				: in std_logic;						-- Input signal
		o_placeholder				: in std_logic;						-- Output signal
	);
end placeholder;

architecture Behavioral of placeholder is
	signal placeholder			: std_logic;

begin

end architecture Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity CPU_random_control_logic_test is
	Port(
		i_clk: in STD_LOGIC;
		i_test_vector: in STD_LOGIC_VECTOR(60 downto 0);
		i_rdy: in STD_LOGIC;
		o_dl_to_db: out STD_LOGIC;
		o_dl_to_adl: out STD_LOGIC;
		o_dl_to_adh: out STD_LOGIC;
		o_O_to_adh0: out STD_LOGIC;
		o_O_to_adh1_7: out STD_LOGIC;
		o_adh_to_abh: out STD_LOGIC;
		o_adl_to_abl: out STD_LOGIC;
		o_pcl_to_pcl: out STD_LOGIC;
		o_adl_to_pcl: out STD_LOGIC;
		o_i_to_pc: out STD_LOGIC;
		o_pcl_to_db: out STD_LOGIC;
		o_pcl_to_adl: out STD_LOGIC;
		o_pch_to_pch: out STD_LOGIC;
		o_adh_to_pch: out STD_LOGIC;
		o_pch_to_db: out STD_LOGIC;
		o_pch_to_adh: out STD_LOGIC;
		o_sb_to_adh: out STD_LOGIC;
		o_sb_to_db: out STD_LOGIC;
		o_O_to_adl0: out STD_LOGIC;
		o_O_to_adl1: out STD_LOGIC;
		o_O_to_adl2: out STD_LOGIC;
		o_s_to_adl: out STD_LOGIC;
		o_sb_to_s: out STD_LOGIC;
		o_s_to_s: out STD_LOGIC;
		o_s_to_sb: out STD_LOGIC;
		o_db_bar_to_add: out STD_LOGIC;
		o_db_to_add: out STD_LOGIC;
		o_adl_to_add: out STD_LOGIC;
		o_i_to_addc: out STD_LOGIC;
		o_sum_select: out STD_LOGIC;
		o_and_select: out STD_LOGIC;
		o_eor_select: out STD_LOGIC;
		o_or_select: out STD_LOGIC;
		o_shift_right_select: out STD_LOGIC;
		o_add_to_adl: out STD_LOGIC;
		o_add_to_sb_0_6: out STD_LOGIC;
		o_add_to_sb_7: out STD_LOGIC;
		o_O_to_add: out STD_LOGIC;
		o_sb_to_add: out STD_LOGIC;
		o_sb_to_ac: out STD_LOGIC;
		o_ac_to_db: out STD_LOGIC;
		o_ac_to_sb: out STD_LOGIC;
		o_sb_to_x: out STD_LOGIC;
		o_x_to_sb: out STD_LOGIC;
		o_sb_to_y: out STD_LOGIC;
		o_y_to_sb: out STD_LOGIC;
		o_p_to_db: out STD_LOGIC;
		o_db0_to_c: out STD_LOGIC;
		o_ir5_to_c: out STD_LOGIC;
		o_acr_to_c: out STD_LOGIC;
		o_db1_to_z: out STD_LOGIC;
		o_dbz_to_z: out STD_LOGIC;
		o_db2_to_i: out STD_LOGIC;
		o_ir5_to_i: out STD_LOGIC;
		o_db3_to_d: out STD_LOGIC;
		o_ir5_to_d: out STD_LOGIC;
		o_db6_to_v: out STD_LOGIC;
		o_avr_to_v: out STD_LOGIC;
		o_i_to_v: out STD_LOGIC;
		o_db7_to_n:out STD_LOGIC;
		o_read_write:out STD_LOGIC);
	end CPU_random_control_logic_test;

architecture Dataflow of CPU_random_control_logic_test is
begin
	o_dl_to_db <= i_test_vector(0);
	o_dl_to_adl <= i_test_vector(1);
	o_dl_to_adh <= i_test_vector(2);
	o_O_to_adh0 <= i_test_vector(3);
	o_O_to_adh1_7 <= i_test_vector(4);
	o_adh_to_abh <= i_test_vector(5);
	o_adl_to_abl <= i_test_vector(6);
	o_pcl_to_pcl <= i_test_vector(7);
	o_adl_to_pcl <= i_test_vector(8);
	o_i_to_pc <= i_test_vector(9);
	o_pcl_to_db <= i_test_vector(10);
	o_pcl_to_adl <= i_test_vector(11);
	o_pch_to_pch <= i_test_vector(12);
	o_adh_to_pch <= i_test_vector(13);
	o_pch_to_db <= i_test_vector(14);
	o_pch_to_adh <= i_test_vector(15);
	o_sb_to_adh <= i_test_vector(16);
	o_sb_to_db <= i_test_vector(17);
	o_O_to_adl0 <= i_test_vector(18);
	o_O_to_adl1 <= i_test_vector(19);
	o_O_to_adl2 <= i_test_vector(20);
	o_s_to_adl <= i_test_vector(21);
	o_sb_to_s <= i_test_vector(22);
	o_s_to_s <= i_test_vector(23);
	o_s_to_sb <= i_test_vector(24);
	o_db_bar_to_add <= i_test_vector(25);
	o_db_to_add <= i_test_vector(26);
	o_adl_to_add <= i_test_vector(27);
	o_i_to_addc <= i_test_vector(28);
	o_sum_select <= i_test_vector(29);
	o_and_select <= i_test_vector(30);
	o_eor_select <= i_test_vector(31);
	o_or_select <= i_test_vector(32);
	o_shift_right_select <= i_test_vector(33);
	o_add_to_adl <= i_test_vector(34);
	o_add_to_sb_0_6 <= i_test_vector(35);
	o_add_to_sb_7 <= i_test_vector(36);
	o_O_to_add <= i_test_vector(37);
	o_sb_to_add <= i_test_vector(38);
	o_sb_to_ac <= i_test_vector(39);
	o_ac_to_db <= i_test_vector(40);
	o_ac_to_sb <= i_test_vector(41);
	o_sb_to_x <= i_test_vector(42);
	o_x_to_sb <= i_test_vector(43);
	o_sb_to_y <= i_test_vector(44);
	o_y_to_sb <= i_test_vector(45);
	o_p_to_db <= i_test_vector(46);
	o_db0_to_c <= i_test_vector(47);
	o_ir5_to_c <= i_test_vector(48);
	o_acr_to_c <= i_test_vector(49);
	o_db1_to_z <= i_test_vector(50);
	o_dbz_to_z <= i_test_vector(51);
	o_db2_to_i <= i_test_vector(52);
	o_ir5_to_i <= i_test_vector(53);
	o_db3_to_d <= i_test_vector(54);
	o_ir5_to_d <= i_test_vector(55);
	o_db6_to_v <= i_test_vector(56);
	o_avr_to_v <= i_test_vector(57);
	o_i_to_v <= i_test_vector(58);
	o_db7_to_n <= i_test_vector(59);
	o_read_write <= i_test_vector(60);
	end Dataflow;
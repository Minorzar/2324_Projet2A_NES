library ieee ;
use ieee.std_logic_1164.all ;
use ieee.numeric_std.all ;

entity CPU_random_control_logic_tb is
end CPU_random_control_logic_tb ;

architecture testbench of CPU_random_control_logic_tb is

	component CPU_random_control_logic
		port(
		
			i_clk							: in std_logic ;
			i_rdy							: in std_logic ;
			i_phi1						: in std_logic ;
			i_phi2						: in std_logic ;
			i_set_overflow				: in std_logic ;
			i_dr							: in unsigned(129 downto 0) ; --the decode ROM array
			i_reset						: in std_logic ;
			i_reset_in_progress		: in std_logic ;
			i_break_in_progress		: in std_logic ;
			i_implied_addressing		: in std_logic ;
			i_two_cycle					: in std_logic ;
			i_t0							: in std_logic ;
			i_ir5							: in std_logic ;
			i_db7							: in std_logic ;
			i_alu_carry_out			: in std_logic ;
			i_break_done				: in std_logic ;
			i_zero_adl0					: in std_logic ;
			i_p_register				: in std_logic_vector(7 downto 0) ;
			o_dl_to_db					: out std_logic ;
			o_dl_to_adl					: out std_logic ;
			o_dl_to_adh					: out std_logic ;
			o_O_to_adh0					: out std_logic ;
			o_O_to_adh1_7				: out std_logic ;
			o_adh_to_abh				: out std_logic ;
			o_adl_to_abl				: out std_logic ;
			o_pcl_to_pcl				: out std_logic ;
			o_adl_to_pcl				: out std_logic ;
			o_i_to_pc					: out std_logic ;
			o_pcl_to_db					: out std_logic ;
			o_pcl_to_adl				: out std_logic ;
			o_pch_to_pch				: out std_logic ;
			o_adh_to_pch				: out std_logic ;
			b_pch_to_db					: buffer std_logic ;
			o_pch_to_adh				: out std_logic ;
			o_sb_to_adh					: out std_logic ;
			o_sb_to_db					: out std_logic ;
			o_O_to_adl0					: out std_logic ;
			o_O_to_adl1					: out std_logic ;
			o_O_to_adl2					: out std_logic ;
			o_s_to_adl					: out std_logic ;
			o_sb_to_s					: out std_logic ;
			o_s_to_s						: out std_logic ;
			o_s_to_sb					: out std_logic ;
			o_db_bar_to_add			: out std_logic ;
			o_db_to_add					: out std_logic ;
			o_adl_to_add				: out std_logic ;
			o_i_to_addc					: out std_logic ;
			o_sum_select				: out std_logic ;
			o_and_select				: out std_logic ;
			o_eor_select				: out std_logic ;
			o_or_select					: out std_logic ;
			o_shift_right_select		: out std_logic ;
			o_add_to_adl				: out std_logic ;
			o_add_to_sb_0_6			: out std_logic ;
			o_add_to_sb_7				: out std_logic ;
			o_O_to_add					: out std_logic ;
			o_sb_to_add					: out std_logic ;
			o_sb_to_ac					: out std_logic ;
			o_ac_to_db					: out std_logic ;
			o_ac_to_sb					: out std_logic ;
			o_sb_to_x					: out std_logic ;
			o_x_to_sb					: out std_logic ;
			o_sb_to_y					: out std_logic ;
			o_y_to_sb					: out std_logic ;
			o_p_to_db					: out std_logic ;
			o_db0_to_c					: out std_logic ;
			o_ir5_to_c					: out std_logic ;
			b_acr_to_c					: buffer std_logic ;
			o_db1_to_z					: out std_logic ;
			b_dbz_to_z					: buffer std_logic ;
			o_db2_to_i					: out std_logic ;
			o_ir5_to_i					: out std_logic ;
			o_db3_to_d					: out std_logic ;
			o_ir5_to_d					: out std_logic ;
			o_db6_to_v					: out std_logic ;
			o_avr_to_v					: out std_logic ;
			o_0_to_v						: out std_logic ;
			o_1_to_v						: out std_logic ;
			o_i_to_v						: out std_logic ;
			o_db7_to_n					: out std_logic ;
			b_t1_reset					: buffer std_logic ;
			o_read_write				: out std_logic
			
		) ;
		
	end component ;
	
	constant clk_period : time := 500ns ;
	
	signal Si_clk: std_logic ;
	signal Si_rdy: std_logic ;
	signal Si_phi1: std_logic ;
	signal Si_phi2: std_logic ;
	signal Si_set_overflow: std_logic ;
	signal Si_dr: unsigned(129 downto 0) ;
	signal Si_reset: std_logic ;
	signal Si_reset_in_progress:  std_logic ;
	signal Si_break_in_progress:  std_logic ;
	signal Si_implied_addressing:  std_logic ;
	signal Si_two_cycle: std_logic ;
	signal Si_t0: std_logic ;
	signal Si_ir5: std_logic ;
	signal Si_db7: std_logic ;
	signal Si_alu_carry_out: std_logic ;
	signal Si_break_done: std_logic ;
	signal Si_zero_adl0: std_logic ;
	signal Si_p_register: std_logic_vector(7 downto 0) ;
	signal So_dl_to_db: std_logic ;
	signal So_dl_to_adl: std_logic ;
	signal So_dl_to_adh: std_logic ;
	signal So_O_to_adh0: std_logic ;
	signal So_O_to_adh1_7: std_logic ;
	signal So_adh_to_abh: std_logic ;
	signal So_adl_to_abl: std_logic ;
	signal So_pcl_to_pcl: std_logic ;
	signal So_adl_to_pcl: std_logic ;
	signal So_i_to_pc: std_logic ;
	signal So_pcl_to_db: std_logic ;
	signal So_pcl_to_adl: std_logic ;
	signal So_pch_to_pch: std_logic ;
	signal So_adh_to_pch: std_logic ;
	signal Sb_pch_to_db: std_logic ;
	signal So_pch_to_adh: std_logic ;
	signal So_sb_to_adh: std_logic ;
	signal So_sb_to_db: std_logic ;
	signal So_O_to_adl0: std_logic ;
	signal So_O_to_adl1: std_logic ;
	signal So_O_to_adl2: std_logic ;
	signal So_s_to_adl: std_logic ;
	signal So_sb_to_s: std_logic ;
	signal So_s_to_s: std_logic ;
	signal So_s_to_sb: std_logic ;
	signal So_db_bar_to_add: std_logic ;
	signal So_db_to_add: std_logic ;
	signal So_adl_to_add: std_logic ;
	signal So_i_to_addc: std_logic ;
	signal So_sum_select: std_logic ;
	signal So_and_select: std_logic ;
	signal So_eor_select: std_logic ;
	signal So_or_select: std_logic ;
	signal So_shift_right_select: std_logic ;
	signal So_add_to_adl: std_logic ;
	signal So_add_to_sb_0_6: std_logic ;
	signal So_add_to_sb_7: std_logic ;
	signal So_O_to_add: std_logic ;
	signal So_sb_to_add: std_logic ;
	signal So_sb_to_ac: std_logic ;
	signal So_ac_to_db: std_logic ;
	signal So_ac_to_sb: std_logic ;
	signal So_sb_to_x: std_logic ;
	signal So_x_to_sb: std_logic ;
	signal So_sb_to_y: std_logic ;
	signal So_y_to_sb: std_logic ;
	signal So_p_to_db: std_logic ;
	signal So_db0_to_c: std_logic ;
	signal So_ir5_to_c: std_logic ;
	signal Sb_acr_to_c: std_logic ;
	signal So_db1_to_z: std_logic ;
	signal Sb_dbz_to_z: std_logic ;
	signal So_db2_to_i: std_logic ;
	signal So_ir5_to_i: std_logic ;
	signal So_db3_to_d: std_logic ;
	signal So_ir5_to_d: std_logic ;
	signal So_db6_to_v: std_logic ;
	signal So_avr_to_v: std_logic ;
	signal So_0_to_v: std_logic ;
	signal So_1_to_v: std_logic ;
	signal So_i_to_v: std_logic ;
	signal So_db7_to_n:std_logic ;
	signal Sb_t1_reset:std_logic ;
	signal So_read_write:std_logic ;
	
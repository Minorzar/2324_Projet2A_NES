library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all; 

entity serialiser_tb is
end serialiser_tb; 

constant CLK_PERIOD : time :=5 ns
signal finished : boolean :=false;



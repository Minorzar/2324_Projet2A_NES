-- ready_control.vhd
--
-- This VHDL module implements "Ready Control".
--
-- Description:
--	

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ready_control is
	Port (
		i_placeholder				: in std_logic;						-- Input signal
		o_placeholder				: in std_logic;						-- Output signal
	);
end ready_control;

architecture Behavioral of ready_control is
	signal placeholder			: std_logic;
begin

end Behavioral;
